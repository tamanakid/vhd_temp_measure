-- pack_temp_conv.vhd
-- package to provide functions, procedures and data types for temperature conversion 



library ieee;
use ieee.std_logic_1164.all;



package pack_temp_conv is
  
  -- temperature units
  type t_unit is (celsius, kelvin, fahrenheit);
  
end package;
